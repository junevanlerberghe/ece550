module register_32(enable, data, result);
	input enable;
	input [31:0] data;
	
	input [31:0] result;